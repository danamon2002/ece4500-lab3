library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity toplevel is
	port( -- TODO: ADD INPUTS AND OUTPUTS
	     );
end entity toplevel;


architecture top of toplevel is

begin



end toplevel;